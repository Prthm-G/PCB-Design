CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 0 30 100 9
0 71 2560 1032
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
62 C:\Users\Manu_\OneDrive\Elec_301\CircuitMaker60S\CM60S\BOM.DAT
0 7
0 71 2560 1032
211288083 384
0
6 Title:
5 Name:
0
0
0
10
7 Ground~
168 333 360 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
12 NPN Trans:B~
219 567 279 0 3 7
0 5 3 2
0
0 0 848 512
6 2N3904
-64 0 -22 8
2 Q2
-50 -10 -36 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
4441 0 0
0
0
12 NPN Trans:B~
219 373 279 0 3 7
0 4 6 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3618 0 0
0
0
10 Capacitor~
219 495 207 0 2 5
0 5 6
0
0 0 848 180
4 22nF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 432 171 0 2 5
0 3 4
0
0 0 848 180
4 22nF
-14 -18 14 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
9 V Source~
197 135 162 0 2 5
0 7 2
0
0 0 17264 0
3 12V
13 0 34 8
2 P1
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
7734 0 0
0
0
9 Resistor~
219 675 90 0 2 5
0 7 3
0
0 0 880 270
4 100k
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 558 90 0 2 5
0 5 7
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 378 90 0 2 5
0 4 7
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 243 90 0 2 5
0 6 7
0
0 0 880 90
4 100k
1 0 29 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
15
1 0 2 0 0 4096 0 1 0 0 12 2
333 354
333 315
1 0 3 0 0 4224 0 5 0 0 15 2
441 171
675 171
2 0 4 0 0 4096 0 5 0 0 13 2
423 171
378 171
1 0 5 0 0 4096 0 4 0 0 6 2
504 207
558 207
2 0 6 0 0 4224 0 4 0 0 14 4
486 207
248 207
248 208
243 208
1 1 5 0 0 4224 0 2 8 0 0 2
558 261
558 108
2 0 7 0 0 4096 0 8 0 0 10 2
558 72
558 46
2 0 7 0 0 0 0 9 0 0 10 2
378 72
378 46
2 0 7 0 0 0 0 10 0 0 10 2
243 72
243 46
1 1 7 0 0 8320 0 6 7 0 0 4
135 141
135 46
675 46
675 72
3 0 2 0 0 0 0 3 0 0 12 2
378 297
378 315
3 2 2 0 0 8320 0 2 6 0 0 4
558 297
558 315
135 315
135 183
1 1 4 0 0 4224 0 9 3 0 0 2
378 108
378 261
2 1 6 0 0 0 0 3 10 0 0 3
355 279
243 279
243 108
2 2 3 0 0 0 0 7 2 0 0 3
675 108
675 279
581 279
0
0
21 0 1
0
0
2 P1
0 5 0.1
0
0 0 0
10 1 1 100000
0 0.05 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
594120 1210432 100 100 0 0
0 0 0 0
68 76 229 146
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
0
1116144 8550464 100 100 0 0
77 66 2507 876
0 71 2560 1032
2507 66
77 66
2507 72
2507 553
0 0
0.05 0 17.88 7.2 0.05 0.05
12393 0
4 1e-006 10
1
558 177
0 5 0 0 1	0 6 0 0
397168 2259008 100 100 0 0
77 66 587 216
640 375 1280 679
587 66
77 66
587 66
587 216
0 0
5 0 1 -0.2 5 5
12401 0
4 1 2
3
378 221
0 4 0 0 1	0 13 0 0
558 238
0 5 0 0 1	0 6 0 0
675 260
0 3 0 0 1	0 15 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
